-- system.vhd

-- Generated using ACDS version 15.0 153

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system is
	port (
		camera_controller_current_frame     : out   std_logic_vector(31 downto 0);                    --       camera_controller.current_frame
		camera_controller_read_done         : in    std_logic                     := '0';             --                        .read_done
		camera_input_clk                    : in    std_logic                     := '0';             --            camera_input.clk
		camera_input_frame_valid            : in    std_logic                     := '0';             --                        .frame_valid
		camera_input_line_valid             : in    std_logic                     := '0';             --                        .line_valid
		camera_input_data                   : in    std_logic_vector(11 downto 0) := (others => '0'); --                        .data
		camera_input_cam_reset_n            : out   std_logic;                                        --                        .cam_reset_n
		clk_clk                             : in    std_logic                     := '0';             --                     clk.clk
		frame_rdy_irq                       : out   std_logic;                                        --               frame_rdy.irq
		i2c_scl                             : inout std_logic                     := '0';             --                     i2c.scl
		i2c_sda                             : inout std_logic                     := '0';             --                        .sda
		sdram_clk_clk                       : out   std_logic;                                        --               sdram_clk.clk
		sdram_wire_addr                     : out   std_logic_vector(12 downto 0);                    --              sdram_wire.addr
		sdram_wire_ba                       : out   std_logic_vector(1 downto 0);                     --                        .ba
		sdram_wire_cas_n                    : out   std_logic;                                        --                        .cas_n
		sdram_wire_cke                      : out   std_logic;                                        --                        .cke
		sdram_wire_cs_n                     : out   std_logic;                                        --                        .cs_n
		sdram_wire_dq                       : inout std_logic_vector(15 downto 0) := (others => '0'); --                        .dq
		sdram_wire_dqm                      : out   std_logic_vector(1 downto 0);                     --                        .dqm
		sdram_wire_ras_n                    : out   std_logic;                                        --                        .ras_n
		sdram_wire_we_n                     : out   std_logic;                                        --                        .we_n
		sensor_output_generator_frame_valid : out   std_logic;                                        -- sensor_output_generator.frame_valid
		sensor_output_generator_line_valid  : out   std_logic;                                        --                        .line_valid
		sensor_output_generator_data        : out   std_logic_vector(11 downto 0)                     --                        .data
	);
end entity system;

architecture rtl of system is
	component CameraController is
		port (
			Clk              : in  std_logic                     := 'X';             -- clk
			AS_Address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			AS_ChipSelect    : in  std_logic                     := 'X';             -- chipselect
			AS_Read          : in  std_logic                     := 'X';             -- read
			AS_Write         : in  std_logic                     := 'X';             -- write
			AS_ReadData      : out std_logic_vector(31 downto 0);                    -- readdata
			AS_WriteData     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nReset           : in  std_logic                     := 'X';             -- reset_n
			CurrentFrame     : out std_logic_vector(31 downto 0);                    -- current_frame
			ReadDone         : in  std_logic                     := 'X';             -- read_done
			AM_Address       : out std_logic_vector(31 downto 0);                    -- address
			AM_ByteEnable    : out std_logic_vector(1 downto 0);                     -- byteenable
			AM_Write         : out std_logic;                                        -- write
			AM_Read          : out std_logic;                                        -- read
			AM_DataWrite     : out std_logic_vector(15 downto 0);                    -- writedata
			AM_DataRead      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			AM_WaitRequest   : in  std_logic                     := 'X';             -- waitrequest
			AM_BurstCount    : out std_logic_vector(2 downto 0);                     -- burstcount
			AM_ReadDataValid : in  std_logic                     := 'X';             -- readdatavalid
			FrameRDY         : out std_logic;                                        -- irq
			CamClk           : in  std_logic                     := 'X';             -- clk
			CamFV            : in  std_logic                     := 'X';             -- frame_valid
			CamLV            : in  std_logic                     := 'X';             -- line_valid
			CamData          : in  std_logic_vector(11 downto 0) := (others => 'X'); -- data
			CamReset_n       : out std_logic                                         -- cam_reset_n
		);
	end component CameraController;

	component system_clocks is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component system_clocks;

	component cmos_sensor_output_generator is
		generic (
			PIX_DEPTH : positive := 8
		);
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			addr        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read        : in  std_logic                     := 'X';             -- read
			write       : in  std_logic                     := 'X';             -- write
			rddata      : out std_logic_vector(31 downto 0);                    -- readdata
			wrdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			frame_valid : out std_logic;                                        -- frame_valid
			line_valid  : out std_logic;                                        -- line_valid
			data        : out std_logic_vector(11 downto 0)                     -- data
		);
	end component cmos_sensor_output_generator;

	component i2c_interface is
		port (
			clk        : in    std_logic                    := 'X';             -- clk
			reset      : in    std_logic                    := 'X';             -- reset
			address    : in    std_logic_vector(1 downto 0) := (others => 'X'); -- address
			chipselect : in    std_logic                    := 'X';             -- chipselect
			write      : in    std_logic                    := 'X';             -- write
			writedata  : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			read       : in    std_logic                    := 'X';             -- read
			readdata   : out   std_logic_vector(7 downto 0);                    -- readdata
			scl        : inout std_logic                    := 'X';             -- scl
			sda        : inout std_logic                    := 'X';             -- sda
			irq        : out   std_logic                                        -- irq
		);
	end component i2c_interface;

	component system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component system_jtag_uart;

	component system_nios2 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(25 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(25 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component system_nios2;

	component system_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component system_sdram;

	component system_mm_interconnect_0 is
		port (
			clocks_sys_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			camera_controller_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			camera_controller_0_avalon_master_address             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			camera_controller_0_avalon_master_waitrequest         : out std_logic;                                        -- waitrequest
			camera_controller_0_avalon_master_burstcount          : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			camera_controller_0_avalon_master_byteenable          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			camera_controller_0_avalon_master_read                : in  std_logic                     := 'X';             -- read
			camera_controller_0_avalon_master_readdata            : out std_logic_vector(15 downto 0);                    -- readdata
			camera_controller_0_avalon_master_readdatavalid       : out std_logic;                                        -- readdatavalid
			camera_controller_0_avalon_master_write               : in  std_logic                     := 'X';             -- write
			camera_controller_0_avalon_master_writedata           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			nios2_data_master_address                             : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			nios2_data_master_waitrequest                         : out std_logic;                                        -- waitrequest
			nios2_data_master_byteenable                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_data_master_read                                : in  std_logic                     := 'X';             -- read
			nios2_data_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_data_master_write                               : in  std_logic                     := 'X';             -- write
			nios2_data_master_writedata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_data_master_debugaccess                         : in  std_logic                     := 'X';             -- debugaccess
			nios2_instruction_master_address                      : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			nios2_instruction_master_waitrequest                  : out std_logic;                                        -- waitrequest
			nios2_instruction_master_read                         : in  std_logic                     := 'X';             -- read
			nios2_instruction_master_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_instruction_master_readdatavalid                : out std_logic;                                        -- readdatavalid
			camera_controller_0_as_address                        : out std_logic_vector(2 downto 0);                     -- address
			camera_controller_0_as_write                          : out std_logic;                                        -- write
			camera_controller_0_as_read                           : out std_logic;                                        -- read
			camera_controller_0_as_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			camera_controller_0_as_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			camera_controller_0_as_chipselect                     : out std_logic;                                        -- chipselect
			cmos_sensor_output_generator_0_avalon_slave_address   : out std_logic_vector(2 downto 0);                     -- address
			cmos_sensor_output_generator_0_avalon_slave_write     : out std_logic;                                        -- write
			cmos_sensor_output_generator_0_avalon_slave_read      : out std_logic;                                        -- read
			cmos_sensor_output_generator_0_avalon_slave_readdata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cmos_sensor_output_generator_0_avalon_slave_writedata : out std_logic_vector(31 downto 0);                    -- writedata
			i2c_0_avalon_slave_address                            : out std_logic_vector(1 downto 0);                     -- address
			i2c_0_avalon_slave_write                              : out std_logic;                                        -- write
			i2c_0_avalon_slave_read                               : out std_logic;                                        -- read
			i2c_0_avalon_slave_readdata                           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_0_avalon_slave_writedata                          : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_0_avalon_slave_chipselect                         : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                     : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                      : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                : out std_logic;                                        -- chipselect
			nios2_jtag_debug_module_address                       : out std_logic_vector(8 downto 0);                     -- address
			nios2_jtag_debug_module_write                         : out std_logic;                                        -- write
			nios2_jtag_debug_module_read                          : out std_logic;                                        -- read
			nios2_jtag_debug_module_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_jtag_debug_module_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_jtag_debug_module_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_jtag_debug_module_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			nios2_jtag_debug_module_debugaccess                   : out std_logic;                                        -- debugaccess
			sdram_s1_address                                      : out std_logic_vector(23 downto 0);                    -- address
			sdram_s1_write                                        : out std_logic;                                        -- write
			sdram_s1_read                                         : out std_logic;                                        -- read
			sdram_s1_readdata                                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                    : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                                   : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                   : out std_logic                                         -- chipselect
		);
	end component system_mm_interconnect_0;

	component system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper;

	component system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component system_rst_controller;

	component system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component system_rst_controller_001;

	signal clocks_sys_clk_clk                                                      : std_logic;                     -- clocks:sys_clk_clk -> [camera_controller_0:Clk, cmos_sensor_output_generator_0:clk, i2c_0:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:clocks_sys_clk_clk, nios2:clk, rst_controller:clk, sdram:clk]
	signal nios2_jtag_debug_module_reset_reset                                     : std_logic;                     -- nios2:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	signal camera_controller_0_avalon_master_readdata                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:camera_controller_0_avalon_master_readdata -> camera_controller_0:AM_DataRead
	signal camera_controller_0_avalon_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:camera_controller_0_avalon_master_waitrequest -> camera_controller_0:AM_WaitRequest
	signal camera_controller_0_avalon_master_address                               : std_logic_vector(31 downto 0); -- camera_controller_0:AM_Address -> mm_interconnect_0:camera_controller_0_avalon_master_address
	signal camera_controller_0_avalon_master_byteenable                            : std_logic_vector(1 downto 0);  -- camera_controller_0:AM_ByteEnable -> mm_interconnect_0:camera_controller_0_avalon_master_byteenable
	signal camera_controller_0_avalon_master_read                                  : std_logic;                     -- camera_controller_0:AM_Read -> mm_interconnect_0:camera_controller_0_avalon_master_read
	signal camera_controller_0_avalon_master_readdatavalid                         : std_logic;                     -- mm_interconnect_0:camera_controller_0_avalon_master_readdatavalid -> camera_controller_0:AM_ReadDataValid
	signal camera_controller_0_avalon_master_write                                 : std_logic;                     -- camera_controller_0:AM_Write -> mm_interconnect_0:camera_controller_0_avalon_master_write
	signal camera_controller_0_avalon_master_writedata                             : std_logic_vector(15 downto 0); -- camera_controller_0:AM_DataWrite -> mm_interconnect_0:camera_controller_0_avalon_master_writedata
	signal camera_controller_0_avalon_master_burstcount                            : std_logic_vector(2 downto 0);  -- camera_controller_0:AM_BurstCount -> mm_interconnect_0:camera_controller_0_avalon_master_burstcount
	signal nios2_data_master_readdata                                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	signal nios2_data_master_waitrequest                                           : std_logic;                     -- mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	signal nios2_data_master_debugaccess                                           : std_logic;                     -- nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	signal nios2_data_master_address                                               : std_logic_vector(25 downto 0); -- nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	signal nios2_data_master_byteenable                                            : std_logic_vector(3 downto 0);  -- nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	signal nios2_data_master_read                                                  : std_logic;                     -- nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	signal nios2_data_master_write                                                 : std_logic;                     -- nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	signal nios2_data_master_writedata                                             : std_logic_vector(31 downto 0); -- nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	signal nios2_instruction_master_readdata                                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	signal nios2_instruction_master_waitrequest                                    : std_logic;                     -- mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	signal nios2_instruction_master_address                                        : std_logic_vector(25 downto 0); -- nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	signal nios2_instruction_master_read                                           : std_logic;                     -- nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	signal nios2_instruction_master_readdatavalid                                  : std_logic;                     -- mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	signal mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_readdata  : std_logic_vector(31 downto 0); -- cmos_sensor_output_generator_0:rddata -> mm_interconnect_0:cmos_sensor_output_generator_0_avalon_slave_readdata
	signal mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_address   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:cmos_sensor_output_generator_0_avalon_slave_address -> cmos_sensor_output_generator_0:addr
	signal mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_read      : std_logic;                     -- mm_interconnect_0:cmos_sensor_output_generator_0_avalon_slave_read -> cmos_sensor_output_generator_0:read
	signal mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_write     : std_logic;                     -- mm_interconnect_0:cmos_sensor_output_generator_0_avalon_slave_write -> cmos_sensor_output_generator_0:write
	signal mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_writedata : std_logic_vector(31 downto 0); -- mm_interconnect_0:cmos_sensor_output_generator_0_avalon_slave_writedata -> cmos_sensor_output_generator_0:wrdata
	signal mm_interconnect_0_sdram_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                     : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                  : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                      : std_logic_vector(23 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                         : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                                : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                        : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_camera_controller_0_as_chipselect                     : std_logic;                     -- mm_interconnect_0:camera_controller_0_as_chipselect -> camera_controller_0:AS_ChipSelect
	signal mm_interconnect_0_camera_controller_0_as_readdata                       : std_logic_vector(31 downto 0); -- camera_controller_0:AS_ReadData -> mm_interconnect_0:camera_controller_0_as_readdata
	signal mm_interconnect_0_camera_controller_0_as_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:camera_controller_0_as_address -> camera_controller_0:AS_Address
	signal mm_interconnect_0_camera_controller_0_as_read                           : std_logic;                     -- mm_interconnect_0:camera_controller_0_as_read -> camera_controller_0:AS_Read
	signal mm_interconnect_0_camera_controller_0_as_write                          : std_logic;                     -- mm_interconnect_0:camera_controller_0_as_write -> camera_controller_0:AS_Write
	signal mm_interconnect_0_camera_controller_0_as_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:camera_controller_0_as_writedata -> camera_controller_0:AS_WriteData
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect                : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                  : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest               : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                   : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                     : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_i2c_0_avalon_slave_chipselect                         : std_logic;                     -- mm_interconnect_0:i2c_0_avalon_slave_chipselect -> i2c_0:chipselect
	signal mm_interconnect_0_i2c_0_avalon_slave_readdata                           : std_logic_vector(7 downto 0);  -- i2c_0:readdata -> mm_interconnect_0:i2c_0_avalon_slave_readdata
	signal mm_interconnect_0_i2c_0_avalon_slave_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:i2c_0_avalon_slave_address -> i2c_0:address
	signal mm_interconnect_0_i2c_0_avalon_slave_read                               : std_logic;                     -- mm_interconnect_0:i2c_0_avalon_slave_read -> i2c_0:read
	signal mm_interconnect_0_i2c_0_avalon_slave_write                              : std_logic;                     -- mm_interconnect_0:i2c_0_avalon_slave_write -> i2c_0:write
	signal mm_interconnect_0_i2c_0_avalon_slave_writedata                          : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_0_avalon_slave_writedata -> i2c_0:writedata
	signal mm_interconnect_0_nios2_jtag_debug_module_readdata                      : std_logic_vector(31 downto 0); -- nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	signal mm_interconnect_0_nios2_jtag_debug_module_waitrequest                   : std_logic;                     -- nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios2_jtag_debug_module_debugaccess                   : std_logic;                     -- mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios2_jtag_debug_module_address                       : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	signal mm_interconnect_0_nios2_jtag_debug_module_read                          : std_logic;                     -- mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	signal mm_interconnect_0_nios2_jtag_debug_module_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	signal mm_interconnect_0_nios2_jtag_debug_module_write                         : std_logic;                     -- mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	signal mm_interconnect_0_nios2_jtag_debug_module_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	signal irq_mapper_receiver0_irq                                                : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal nios2_d_irq_irq                                                         : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2:d_irq
	signal rst_controller_reset_out_reset                                          : std_logic;                     -- rst_controller:reset_out -> [cmos_sensor_output_generator_0:reset, i2c_0:reset, irq_mapper:reset, mm_interconnect_0:camera_controller_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                      : std_logic;                     -- rst_controller:reset_req -> [nios2:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                                      : std_logic;                     -- rst_controller_001:reset_out -> clocks:ref_reset_reset
	signal mm_interconnect_0_sdram_s1_read_ports_inv                               : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv            : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv           : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                                : std_logic;                     -- rst_controller_reset_out_reset:inv -> [camera_controller_0:nReset, jtag_uart:rst_n, nios2:reset_n, sdram:reset_n]

begin

	camera_controller_0 : component CameraController
		port map (
			Clk              => clocks_sys_clk_clk,                                  --            clock.clk
			AS_Address       => mm_interconnect_0_camera_controller_0_as_address,    --               as.address
			AS_ChipSelect    => mm_interconnect_0_camera_controller_0_as_chipselect, --                 .chipselect
			AS_Read          => mm_interconnect_0_camera_controller_0_as_read,       --                 .read
			AS_Write         => mm_interconnect_0_camera_controller_0_as_write,      --                 .write
			AS_ReadData      => mm_interconnect_0_camera_controller_0_as_readdata,   --                 .readdata
			AS_WriteData     => mm_interconnect_0_camera_controller_0_as_writedata,  --                 .writedata
			nReset           => rst_controller_reset_out_reset_ports_inv,            --            reset.reset_n
			CurrentFrame     => camera_controller_current_frame,                     --      conduit_end.current_frame
			ReadDone         => camera_controller_read_done,                         --                 .read_done
			AM_Address       => camera_controller_0_avalon_master_address,           --    avalon_master.address
			AM_ByteEnable    => camera_controller_0_avalon_master_byteenable,        --                 .byteenable
			AM_Write         => camera_controller_0_avalon_master_write,             --                 .write
			AM_Read          => camera_controller_0_avalon_master_read,              --                 .read
			AM_DataWrite     => camera_controller_0_avalon_master_writedata,         --                 .writedata
			AM_DataRead      => camera_controller_0_avalon_master_readdata,          --                 .readdata
			AM_WaitRequest   => camera_controller_0_avalon_master_waitrequest,       --                 .waitrequest
			AM_BurstCount    => camera_controller_0_avalon_master_burstcount,        --                 .burstcount
			AM_ReadDataValid => camera_controller_0_avalon_master_readdatavalid,     --                 .readdatavalid
			FrameRDY         => frame_rdy_irq,                                       -- interrupt_sender.irq
			CamClk           => camera_input_clk,                                    --     camera_input.clk
			CamFV            => camera_input_frame_valid,                            --                 .frame_valid
			CamLV            => camera_input_line_valid,                             --                 .line_valid
			CamData          => camera_input_data,                                   --                 .data
			CamReset_n       => camera_input_cam_reset_n                             --                 .cam_reset_n
		);

	clocks : component system_clocks
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => rst_controller_001_reset_out_reset, --    ref_reset.reset
			sys_clk_clk        => clocks_sys_clk_clk,                 --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                      --    sdram_clk.clk
			reset_source_reset => open                                -- reset_source.reset
		);

	cmos_sensor_output_generator_0 : component cmos_sensor_output_generator
		generic map (
			PIX_DEPTH => 12
		)
		port map (
			clk         => clocks_sys_clk_clk,                                                      --        clock.clk
			reset       => rst_controller_reset_out_reset,                                          --        reset.reset
			addr        => mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_address,   -- avalon_slave.address
			read        => mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_read,      --             .read
			write       => mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_write,     --             .write
			rddata      => mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_readdata,  --             .readdata
			wrdata      => mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_writedata, --             .writedata
			frame_valid => sensor_output_generator_frame_valid,                                     --  cmos_sensor.frame_valid
			line_valid  => sensor_output_generator_line_valid,                                      --             .line_valid
			data        => sensor_output_generator_data                                             --             .data
		);

	i2c_0 : component i2c_interface
		port map (
			clk        => clocks_sys_clk_clk,                              --            clock.clk
			reset      => rst_controller_reset_out_reset,                  --            reset.reset
			address    => mm_interconnect_0_i2c_0_avalon_slave_address,    --     avalon_slave.address
			chipselect => mm_interconnect_0_i2c_0_avalon_slave_chipselect, --                 .chipselect
			write      => mm_interconnect_0_i2c_0_avalon_slave_write,      --                 .write
			writedata  => mm_interconnect_0_i2c_0_avalon_slave_writedata,  --                 .writedata
			read       => mm_interconnect_0_i2c_0_avalon_slave_read,       --                 .read
			readdata   => mm_interconnect_0_i2c_0_avalon_slave_readdata,   --                 .readdata
			scl        => i2c_scl,                                         --              i2c.scl
			sda        => i2c_sda,                                         --                 .sda
			irq        => open                                             -- interrupt_sender.irq
		);

	jtag_uart : component system_jtag_uart
		port map (
			clk            => clocks_sys_clk_clk,                                            --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	nios2 : component system_nios2
		port map (
			clk                                   => clocks_sys_clk_clk,                                    --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,              --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                    --                          .reset_req
			d_address                             => nios2_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_data_master_read,                                --                          .read
			d_readdata                            => nios2_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_data_master_write,                               --                          .write
			d_writedata                           => nios2_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_instruction_master_waitrequest,                  --                          .waitrequest
			i_readdatavalid                       => nios2_instruction_master_readdatavalid,                --                          .readdatavalid
			d_irq                                 => nios2_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios2_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios2_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios2_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios2_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios2_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios2_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios2_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios2_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                   -- custom_instruction_master.readra
		);

	sdram : component system_sdram
		port map (
			clk            => clocks_sys_clk_clk,                              --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	mm_interconnect_0 : component system_mm_interconnect_0
		port map (
			clocks_sys_clk_clk                                    => clocks_sys_clk_clk,                                                      --                                  clocks_sys_clk.clk
			camera_controller_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                          -- camera_controller_0_reset_reset_bridge_in_reset.reset
			camera_controller_0_avalon_master_address             => camera_controller_0_avalon_master_address,                               --               camera_controller_0_avalon_master.address
			camera_controller_0_avalon_master_waitrequest         => camera_controller_0_avalon_master_waitrequest,                           --                                                .waitrequest
			camera_controller_0_avalon_master_burstcount          => camera_controller_0_avalon_master_burstcount,                            --                                                .burstcount
			camera_controller_0_avalon_master_byteenable          => camera_controller_0_avalon_master_byteenable,                            --                                                .byteenable
			camera_controller_0_avalon_master_read                => camera_controller_0_avalon_master_read,                                  --                                                .read
			camera_controller_0_avalon_master_readdata            => camera_controller_0_avalon_master_readdata,                              --                                                .readdata
			camera_controller_0_avalon_master_readdatavalid       => camera_controller_0_avalon_master_readdatavalid,                         --                                                .readdatavalid
			camera_controller_0_avalon_master_write               => camera_controller_0_avalon_master_write,                                 --                                                .write
			camera_controller_0_avalon_master_writedata           => camera_controller_0_avalon_master_writedata,                             --                                                .writedata
			nios2_data_master_address                             => nios2_data_master_address,                                               --                               nios2_data_master.address
			nios2_data_master_waitrequest                         => nios2_data_master_waitrequest,                                           --                                                .waitrequest
			nios2_data_master_byteenable                          => nios2_data_master_byteenable,                                            --                                                .byteenable
			nios2_data_master_read                                => nios2_data_master_read,                                                  --                                                .read
			nios2_data_master_readdata                            => nios2_data_master_readdata,                                              --                                                .readdata
			nios2_data_master_write                               => nios2_data_master_write,                                                 --                                                .write
			nios2_data_master_writedata                           => nios2_data_master_writedata,                                             --                                                .writedata
			nios2_data_master_debugaccess                         => nios2_data_master_debugaccess,                                           --                                                .debugaccess
			nios2_instruction_master_address                      => nios2_instruction_master_address,                                        --                        nios2_instruction_master.address
			nios2_instruction_master_waitrequest                  => nios2_instruction_master_waitrequest,                                    --                                                .waitrequest
			nios2_instruction_master_read                         => nios2_instruction_master_read,                                           --                                                .read
			nios2_instruction_master_readdata                     => nios2_instruction_master_readdata,                                       --                                                .readdata
			nios2_instruction_master_readdatavalid                => nios2_instruction_master_readdatavalid,                                  --                                                .readdatavalid
			camera_controller_0_as_address                        => mm_interconnect_0_camera_controller_0_as_address,                        --                          camera_controller_0_as.address
			camera_controller_0_as_write                          => mm_interconnect_0_camera_controller_0_as_write,                          --                                                .write
			camera_controller_0_as_read                           => mm_interconnect_0_camera_controller_0_as_read,                           --                                                .read
			camera_controller_0_as_readdata                       => mm_interconnect_0_camera_controller_0_as_readdata,                       --                                                .readdata
			camera_controller_0_as_writedata                      => mm_interconnect_0_camera_controller_0_as_writedata,                      --                                                .writedata
			camera_controller_0_as_chipselect                     => mm_interconnect_0_camera_controller_0_as_chipselect,                     --                                                .chipselect
			cmos_sensor_output_generator_0_avalon_slave_address   => mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_address,   --     cmos_sensor_output_generator_0_avalon_slave.address
			cmos_sensor_output_generator_0_avalon_slave_write     => mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_write,     --                                                .write
			cmos_sensor_output_generator_0_avalon_slave_read      => mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_read,      --                                                .read
			cmos_sensor_output_generator_0_avalon_slave_readdata  => mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_readdata,  --                                                .readdata
			cmos_sensor_output_generator_0_avalon_slave_writedata => mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_writedata, --                                                .writedata
			i2c_0_avalon_slave_address                            => mm_interconnect_0_i2c_0_avalon_slave_address,                            --                              i2c_0_avalon_slave.address
			i2c_0_avalon_slave_write                              => mm_interconnect_0_i2c_0_avalon_slave_write,                              --                                                .write
			i2c_0_avalon_slave_read                               => mm_interconnect_0_i2c_0_avalon_slave_read,                               --                                                .read
			i2c_0_avalon_slave_readdata                           => mm_interconnect_0_i2c_0_avalon_slave_readdata,                           --                                                .readdata
			i2c_0_avalon_slave_writedata                          => mm_interconnect_0_i2c_0_avalon_slave_writedata,                          --                                                .writedata
			i2c_0_avalon_slave_chipselect                         => mm_interconnect_0_i2c_0_avalon_slave_chipselect,                         --                                                .chipselect
			jtag_uart_avalon_jtag_slave_address                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,                   --                     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,                     --                                                .write
			jtag_uart_avalon_jtag_slave_read                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                      --                                                .read
			jtag_uart_avalon_jtag_slave_readdata                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,                  --                                                .readdata
			jtag_uart_avalon_jtag_slave_writedata                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,                 --                                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,               --                                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,                --                                                .chipselect
			nios2_jtag_debug_module_address                       => mm_interconnect_0_nios2_jtag_debug_module_address,                       --                         nios2_jtag_debug_module.address
			nios2_jtag_debug_module_write                         => mm_interconnect_0_nios2_jtag_debug_module_write,                         --                                                .write
			nios2_jtag_debug_module_read                          => mm_interconnect_0_nios2_jtag_debug_module_read,                          --                                                .read
			nios2_jtag_debug_module_readdata                      => mm_interconnect_0_nios2_jtag_debug_module_readdata,                      --                                                .readdata
			nios2_jtag_debug_module_writedata                     => mm_interconnect_0_nios2_jtag_debug_module_writedata,                     --                                                .writedata
			nios2_jtag_debug_module_byteenable                    => mm_interconnect_0_nios2_jtag_debug_module_byteenable,                    --                                                .byteenable
			nios2_jtag_debug_module_waitrequest                   => mm_interconnect_0_nios2_jtag_debug_module_waitrequest,                   --                                                .waitrequest
			nios2_jtag_debug_module_debugaccess                   => mm_interconnect_0_nios2_jtag_debug_module_debugaccess,                   --                                                .debugaccess
			sdram_s1_address                                      => mm_interconnect_0_sdram_s1_address,                                      --                                        sdram_s1.address
			sdram_s1_write                                        => mm_interconnect_0_sdram_s1_write,                                        --                                                .write
			sdram_s1_read                                         => mm_interconnect_0_sdram_s1_read,                                         --                                                .read
			sdram_s1_readdata                                     => mm_interconnect_0_sdram_s1_readdata,                                     --                                                .readdata
			sdram_s1_writedata                                    => mm_interconnect_0_sdram_s1_writedata,                                    --                                                .writedata
			sdram_s1_byteenable                                   => mm_interconnect_0_sdram_s1_byteenable,                                   --                                                .byteenable
			sdram_s1_readdatavalid                                => mm_interconnect_0_sdram_s1_readdatavalid,                                --                                                .readdatavalid
			sdram_s1_waitrequest                                  => mm_interconnect_0_sdram_s1_waitrequest,                                  --                                                .waitrequest
			sdram_s1_chipselect                                   => mm_interconnect_0_sdram_s1_chipselect                                    --                                                .chipselect
		);

	irq_mapper : component system_irq_mapper
		port map (
			clk           => clocks_sys_clk_clk,             --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios2_d_irq_irq                 --    sender.irq
		);

	rst_controller : component system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1      => nios2_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => clocks_sys_clk_clk,                  --       clk.clk
			reset_out      => rst_controller_reset_out_reset,      -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,  --          .reset_req
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_in2      => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	rst_controller_001 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_jtag_debug_module_reset_reset, -- reset_in0.reset
			clk            => clk_clk,                             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                                -- (terminated)
			reset_req_in0  => '0',                                 -- (terminated)
			reset_in1      => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_in2      => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of system
