// system.v

// Generated using ACDS version 15.0 153

`timescale 1 ps / 1 ps
module system (
		output wire [31:0] camera_controller_current_frame,     //       camera_controller.current_frame
		input  wire        camera_controller_read_done,         //                        .read_done
		input  wire        camera_input_clk,                    //            camera_input.clk
		input  wire        camera_input_frame_valid,            //                        .frame_valid
		input  wire        camera_input_line_valid,             //                        .line_valid
		input  wire [11:0] camera_input_data,                   //                        .data
		output wire        camera_input_cam_reset_n,            //                        .cam_reset_n
		input  wire        clk_clk,                             //                     clk.clk
		output wire        frame_rdy_irq,                       //               frame_rdy.irq
		inout  wire        i2c_scl,                             //                     i2c.scl
		inout  wire        i2c_sda,                             //                        .sda
		output wire        sdram_clk_clk,                       //               sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                     //              sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                       //                        .ba
		output wire        sdram_wire_cas_n,                    //                        .cas_n
		output wire        sdram_wire_cke,                      //                        .cke
		output wire        sdram_wire_cs_n,                     //                        .cs_n
		inout  wire [15:0] sdram_wire_dq,                       //                        .dq
		output wire [1:0]  sdram_wire_dqm,                      //                        .dqm
		output wire        sdram_wire_ras_n,                    //                        .ras_n
		output wire        sdram_wire_we_n,                     //                        .we_n
		output wire        sensor_output_generator_frame_valid, // sensor_output_generator.frame_valid
		output wire        sensor_output_generator_line_valid,  //                        .line_valid
		output wire [11:0] sensor_output_generator_data         //                        .data
	);

	wire         clocks_sys_clk_clk;                                                      // clocks:sys_clk_clk -> [camera_controller_0:Clk, cmos_sensor_output_generator_0:clk, i2c_0:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:clocks_sys_clk_clk, nios2:clk, rst_controller:clk, sdram:clk]
	wire         nios2_jtag_debug_module_reset_reset;                                     // nios2:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire  [15:0] camera_controller_0_avalon_master_readdata;                              // mm_interconnect_0:camera_controller_0_avalon_master_readdata -> camera_controller_0:AM_DataRead
	wire         camera_controller_0_avalon_master_waitrequest;                           // mm_interconnect_0:camera_controller_0_avalon_master_waitrequest -> camera_controller_0:AM_WaitRequest
	wire  [31:0] camera_controller_0_avalon_master_address;                               // camera_controller_0:AM_Address -> mm_interconnect_0:camera_controller_0_avalon_master_address
	wire   [1:0] camera_controller_0_avalon_master_byteenable;                            // camera_controller_0:AM_ByteEnable -> mm_interconnect_0:camera_controller_0_avalon_master_byteenable
	wire         camera_controller_0_avalon_master_read;                                  // camera_controller_0:AM_Read -> mm_interconnect_0:camera_controller_0_avalon_master_read
	wire         camera_controller_0_avalon_master_readdatavalid;                         // mm_interconnect_0:camera_controller_0_avalon_master_readdatavalid -> camera_controller_0:AM_ReadDataValid
	wire         camera_controller_0_avalon_master_write;                                 // camera_controller_0:AM_Write -> mm_interconnect_0:camera_controller_0_avalon_master_write
	wire  [15:0] camera_controller_0_avalon_master_writedata;                             // camera_controller_0:AM_DataWrite -> mm_interconnect_0:camera_controller_0_avalon_master_writedata
	wire   [2:0] camera_controller_0_avalon_master_burstcount;                            // camera_controller_0:AM_BurstCount -> mm_interconnect_0:camera_controller_0_avalon_master_burstcount
	wire  [31:0] nios2_data_master_readdata;                                              // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                                           // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                                           // nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [25:0] nios2_data_master_address;                                               // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                            // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                                  // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                                                 // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                             // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                                       // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                                    // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [25:0] nios2_instruction_master_address;                                        // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                           // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire         nios2_instruction_master_readdatavalid;                                  // mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	wire  [31:0] mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_readdata;  // cmos_sensor_output_generator_0:rddata -> mm_interconnect_0:cmos_sensor_output_generator_0_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_address;   // mm_interconnect_0:cmos_sensor_output_generator_0_avalon_slave_address -> cmos_sensor_output_generator_0:addr
	wire         mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_read;      // mm_interconnect_0:cmos_sensor_output_generator_0_avalon_slave_read -> cmos_sensor_output_generator_0:read
	wire         mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_write;     // mm_interconnect_0:cmos_sensor_output_generator_0_avalon_slave_write -> cmos_sensor_output_generator_0:write
	wire  [31:0] mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_writedata; // mm_interconnect_0:cmos_sensor_output_generator_0_avalon_slave_writedata -> cmos_sensor_output_generator_0:wrdata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                   // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                     // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                  // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                                      // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                         // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                   // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                        // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                    // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_camera_controller_0_as_chipselect;                     // mm_interconnect_0:camera_controller_0_as_chipselect -> camera_controller_0:AS_ChipSelect
	wire  [31:0] mm_interconnect_0_camera_controller_0_as_readdata;                       // camera_controller_0:AS_ReadData -> mm_interconnect_0:camera_controller_0_as_readdata
	wire   [2:0] mm_interconnect_0_camera_controller_0_as_address;                        // mm_interconnect_0:camera_controller_0_as_address -> camera_controller_0:AS_Address
	wire         mm_interconnect_0_camera_controller_0_as_read;                           // mm_interconnect_0:camera_controller_0_as_read -> camera_controller_0:AS_Read
	wire         mm_interconnect_0_camera_controller_0_as_write;                          // mm_interconnect_0:camera_controller_0_as_write -> camera_controller_0:AS_Write
	wire  [31:0] mm_interconnect_0_camera_controller_0_as_writedata;                      // mm_interconnect_0:camera_controller_0_as_writedata -> camera_controller_0:AS_WriteData
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                  // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;               // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_i2c_0_avalon_slave_chipselect;                         // mm_interconnect_0:i2c_0_avalon_slave_chipselect -> i2c_0:chipselect
	wire   [7:0] mm_interconnect_0_i2c_0_avalon_slave_readdata;                           // i2c_0:readdata -> mm_interconnect_0:i2c_0_avalon_slave_readdata
	wire   [1:0] mm_interconnect_0_i2c_0_avalon_slave_address;                            // mm_interconnect_0:i2c_0_avalon_slave_address -> i2c_0:address
	wire         mm_interconnect_0_i2c_0_avalon_slave_read;                               // mm_interconnect_0:i2c_0_avalon_slave_read -> i2c_0:read
	wire         mm_interconnect_0_i2c_0_avalon_slave_write;                              // mm_interconnect_0:i2c_0_avalon_slave_write -> i2c_0:write
	wire   [7:0] mm_interconnect_0_i2c_0_avalon_slave_writedata;                          // mm_interconnect_0:i2c_0_avalon_slave_writedata -> i2c_0:writedata
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_readdata;                      // nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_waitrequest;                   // nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_jtag_debug_module_debugaccess;                   // mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_jtag_debug_module_address;                       // mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_jtag_debug_module_read;                          // mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_jtag_debug_module_byteenable;                    // mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_jtag_debug_module_write;                         // mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_writedata;                     // mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	wire         irq_mapper_receiver0_irq;                                                // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_d_irq_irq;                                                         // irq_mapper:sender_irq -> nios2:d_irq
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [camera_controller_0:nReset, cmos_sensor_output_generator_0:reset, i2c_0:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:camera_controller_0_reset_reset_bridge_in_reset_reset, nios2:reset_n, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [nios2:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> clocks:ref_reset_reset

	CameraController camera_controller_0 (
		.Clk              (clocks_sys_clk_clk),                                  //            clock.clk
		.AS_Address       (mm_interconnect_0_camera_controller_0_as_address),    //               as.address
		.AS_ChipSelect    (mm_interconnect_0_camera_controller_0_as_chipselect), //                 .chipselect
		.AS_Read          (mm_interconnect_0_camera_controller_0_as_read),       //                 .read
		.AS_Write         (mm_interconnect_0_camera_controller_0_as_write),      //                 .write
		.AS_ReadData      (mm_interconnect_0_camera_controller_0_as_readdata),   //                 .readdata
		.AS_WriteData     (mm_interconnect_0_camera_controller_0_as_writedata),  //                 .writedata
		.nReset           (~rst_controller_reset_out_reset),                     //            reset.reset_n
		.CurrentFrame     (camera_controller_current_frame),                     //      conduit_end.current_frame
		.ReadDone         (camera_controller_read_done),                         //                 .read_done
		.AM_Address       (camera_controller_0_avalon_master_address),           //    avalon_master.address
		.AM_ByteEnable    (camera_controller_0_avalon_master_byteenable),        //                 .byteenable
		.AM_Write         (camera_controller_0_avalon_master_write),             //                 .write
		.AM_Read          (camera_controller_0_avalon_master_read),              //                 .read
		.AM_DataWrite     (camera_controller_0_avalon_master_writedata),         //                 .writedata
		.AM_DataRead      (camera_controller_0_avalon_master_readdata),          //                 .readdata
		.AM_WaitRequest   (camera_controller_0_avalon_master_waitrequest),       //                 .waitrequest
		.AM_BurstCount    (camera_controller_0_avalon_master_burstcount),        //                 .burstcount
		.AM_ReadDataValid (camera_controller_0_avalon_master_readdatavalid),     //                 .readdatavalid
		.FrameRDY         (frame_rdy_irq),                                       // interrupt_sender.irq
		.CamClk           (camera_input_clk),                                    //     camera_input.clk
		.CamFV            (camera_input_frame_valid),                            //                 .frame_valid
		.CamLV            (camera_input_line_valid),                             //                 .line_valid
		.CamData          (camera_input_data),                                   //                 .data
		.CamReset_n       (camera_input_cam_reset_n)                             //                 .cam_reset_n
	);

	system_clocks clocks (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_001_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (clocks_sys_clk_clk),                 //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset ()                                    // reset_source.reset
	);

	cmos_sensor_output_generator #(
		.PIX_DEPTH (12)
	) cmos_sensor_output_generator_0 (
		.clk         (clocks_sys_clk_clk),                                                      //        clock.clk
		.reset       (rst_controller_reset_out_reset),                                          //        reset.reset
		.addr        (mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_address),   // avalon_slave.address
		.read        (mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_read),      //             .read
		.write       (mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_write),     //             .write
		.rddata      (mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_readdata),  //             .readdata
		.wrdata      (mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_writedata), //             .writedata
		.frame_valid (sensor_output_generator_frame_valid),                                     //  cmos_sensor.frame_valid
		.line_valid  (sensor_output_generator_line_valid),                                      //             .line_valid
		.data        (sensor_output_generator_data)                                             //             .data
	);

	i2c_interface i2c_0 (
		.clk        (clocks_sys_clk_clk),                              //            clock.clk
		.reset      (rst_controller_reset_out_reset),                  //            reset.reset
		.address    (mm_interconnect_0_i2c_0_avalon_slave_address),    //     avalon_slave.address
		.chipselect (mm_interconnect_0_i2c_0_avalon_slave_chipselect), //                 .chipselect
		.write      (mm_interconnect_0_i2c_0_avalon_slave_write),      //                 .write
		.writedata  (mm_interconnect_0_i2c_0_avalon_slave_writedata),  //                 .writedata
		.read       (mm_interconnect_0_i2c_0_avalon_slave_read),       //                 .read
		.readdata   (mm_interconnect_0_i2c_0_avalon_slave_readdata),   //                 .readdata
		.scl        (i2c_scl),                                         //              i2c.scl
		.sda        (i2c_sda),                                         //                 .sda
		.irq        ()                                                 // interrupt_sender.irq
	);

	system_jtag_uart jtag_uart (
		.clk            (clocks_sys_clk_clk),                                        //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	system_nios2 nios2 (
		.clk                                   (clocks_sys_clk_clk),                                    //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (nios2_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_data_master_read),                                //                          .read
		.d_readdata                            (nios2_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_data_master_write),                               //                          .write
		.d_writedata                           (nios2_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	system_sdram sdram (
		.clk            (clocks_sys_clk_clk),                       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.clocks_sys_clk_clk                                    (clocks_sys_clk_clk),                                                      //                                  clocks_sys_clk.clk
		.camera_controller_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                          // camera_controller_0_reset_reset_bridge_in_reset.reset
		.camera_controller_0_avalon_master_address             (camera_controller_0_avalon_master_address),                               //               camera_controller_0_avalon_master.address
		.camera_controller_0_avalon_master_waitrequest         (camera_controller_0_avalon_master_waitrequest),                           //                                                .waitrequest
		.camera_controller_0_avalon_master_burstcount          (camera_controller_0_avalon_master_burstcount),                            //                                                .burstcount
		.camera_controller_0_avalon_master_byteenable          (camera_controller_0_avalon_master_byteenable),                            //                                                .byteenable
		.camera_controller_0_avalon_master_read                (camera_controller_0_avalon_master_read),                                  //                                                .read
		.camera_controller_0_avalon_master_readdata            (camera_controller_0_avalon_master_readdata),                              //                                                .readdata
		.camera_controller_0_avalon_master_readdatavalid       (camera_controller_0_avalon_master_readdatavalid),                         //                                                .readdatavalid
		.camera_controller_0_avalon_master_write               (camera_controller_0_avalon_master_write),                                 //                                                .write
		.camera_controller_0_avalon_master_writedata           (camera_controller_0_avalon_master_writedata),                             //                                                .writedata
		.nios2_data_master_address                             (nios2_data_master_address),                                               //                               nios2_data_master.address
		.nios2_data_master_waitrequest                         (nios2_data_master_waitrequest),                                           //                                                .waitrequest
		.nios2_data_master_byteenable                          (nios2_data_master_byteenable),                                            //                                                .byteenable
		.nios2_data_master_read                                (nios2_data_master_read),                                                  //                                                .read
		.nios2_data_master_readdata                            (nios2_data_master_readdata),                                              //                                                .readdata
		.nios2_data_master_write                               (nios2_data_master_write),                                                 //                                                .write
		.nios2_data_master_writedata                           (nios2_data_master_writedata),                                             //                                                .writedata
		.nios2_data_master_debugaccess                         (nios2_data_master_debugaccess),                                           //                                                .debugaccess
		.nios2_instruction_master_address                      (nios2_instruction_master_address),                                        //                        nios2_instruction_master.address
		.nios2_instruction_master_waitrequest                  (nios2_instruction_master_waitrequest),                                    //                                                .waitrequest
		.nios2_instruction_master_read                         (nios2_instruction_master_read),                                           //                                                .read
		.nios2_instruction_master_readdata                     (nios2_instruction_master_readdata),                                       //                                                .readdata
		.nios2_instruction_master_readdatavalid                (nios2_instruction_master_readdatavalid),                                  //                                                .readdatavalid
		.camera_controller_0_as_address                        (mm_interconnect_0_camera_controller_0_as_address),                        //                          camera_controller_0_as.address
		.camera_controller_0_as_write                          (mm_interconnect_0_camera_controller_0_as_write),                          //                                                .write
		.camera_controller_0_as_read                           (mm_interconnect_0_camera_controller_0_as_read),                           //                                                .read
		.camera_controller_0_as_readdata                       (mm_interconnect_0_camera_controller_0_as_readdata),                       //                                                .readdata
		.camera_controller_0_as_writedata                      (mm_interconnect_0_camera_controller_0_as_writedata),                      //                                                .writedata
		.camera_controller_0_as_chipselect                     (mm_interconnect_0_camera_controller_0_as_chipselect),                     //                                                .chipselect
		.cmos_sensor_output_generator_0_avalon_slave_address   (mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_address),   //     cmos_sensor_output_generator_0_avalon_slave.address
		.cmos_sensor_output_generator_0_avalon_slave_write     (mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_write),     //                                                .write
		.cmos_sensor_output_generator_0_avalon_slave_read      (mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_read),      //                                                .read
		.cmos_sensor_output_generator_0_avalon_slave_readdata  (mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_readdata),  //                                                .readdata
		.cmos_sensor_output_generator_0_avalon_slave_writedata (mm_interconnect_0_cmos_sensor_output_generator_0_avalon_slave_writedata), //                                                .writedata
		.i2c_0_avalon_slave_address                            (mm_interconnect_0_i2c_0_avalon_slave_address),                            //                              i2c_0_avalon_slave.address
		.i2c_0_avalon_slave_write                              (mm_interconnect_0_i2c_0_avalon_slave_write),                              //                                                .write
		.i2c_0_avalon_slave_read                               (mm_interconnect_0_i2c_0_avalon_slave_read),                               //                                                .read
		.i2c_0_avalon_slave_readdata                           (mm_interconnect_0_i2c_0_avalon_slave_readdata),                           //                                                .readdata
		.i2c_0_avalon_slave_writedata                          (mm_interconnect_0_i2c_0_avalon_slave_writedata),                          //                                                .writedata
		.i2c_0_avalon_slave_chipselect                         (mm_interconnect_0_i2c_0_avalon_slave_chipselect),                         //                                                .chipselect
		.jtag_uart_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                   //                     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                     //                                                .write
		.jtag_uart_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                      //                                                .read
		.jtag_uart_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                  //                                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                 //                                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),               //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                //                                                .chipselect
		.nios2_jtag_debug_module_address                       (mm_interconnect_0_nios2_jtag_debug_module_address),                       //                         nios2_jtag_debug_module.address
		.nios2_jtag_debug_module_write                         (mm_interconnect_0_nios2_jtag_debug_module_write),                         //                                                .write
		.nios2_jtag_debug_module_read                          (mm_interconnect_0_nios2_jtag_debug_module_read),                          //                                                .read
		.nios2_jtag_debug_module_readdata                      (mm_interconnect_0_nios2_jtag_debug_module_readdata),                      //                                                .readdata
		.nios2_jtag_debug_module_writedata                     (mm_interconnect_0_nios2_jtag_debug_module_writedata),                     //                                                .writedata
		.nios2_jtag_debug_module_byteenable                    (mm_interconnect_0_nios2_jtag_debug_module_byteenable),                    //                                                .byteenable
		.nios2_jtag_debug_module_waitrequest                   (mm_interconnect_0_nios2_jtag_debug_module_waitrequest),                   //                                                .waitrequest
		.nios2_jtag_debug_module_debugaccess                   (mm_interconnect_0_nios2_jtag_debug_module_debugaccess),                   //                                                .debugaccess
		.sdram_s1_address                                      (mm_interconnect_0_sdram_s1_address),                                      //                                        sdram_s1.address
		.sdram_s1_write                                        (mm_interconnect_0_sdram_s1_write),                                        //                                                .write
		.sdram_s1_read                                         (mm_interconnect_0_sdram_s1_read),                                         //                                                .read
		.sdram_s1_readdata                                     (mm_interconnect_0_sdram_s1_readdata),                                     //                                                .readdata
		.sdram_s1_writedata                                    (mm_interconnect_0_sdram_s1_writedata),                                    //                                                .writedata
		.sdram_s1_byteenable                                   (mm_interconnect_0_sdram_s1_byteenable),                                   //                                                .byteenable
		.sdram_s1_readdatavalid                                (mm_interconnect_0_sdram_s1_readdatavalid),                                //                                                .readdatavalid
		.sdram_s1_waitrequest                                  (mm_interconnect_0_sdram_s1_waitrequest),                                  //                                                .waitrequest
		.sdram_s1_chipselect                                   (mm_interconnect_0_sdram_s1_chipselect)                                    //                                                .chipselect
	);

	system_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clocks_sys_clk_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_jtag_debug_module_reset_reset), // reset_in0.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
